-------------------------------------------------------------
-- Filename:  CRC32_LUT2ab.VHD
-- Authors: 
-- 	from http://www.xilinx.com/support/documentation/sw_manuals/xilinx14_4/xst_v6s6.pdf  p262
--		Alain Zarembowitch / MSS
-- Version: Rev 0
-- Last modified: 12/13/17
-- Inheritance: 	ROM1.vhd 8/24/16
--
-- description:  synthesizable generic dual port ROM containing two tables of 256 CRC32s values each
-- (called LUT2a and LUT2b)
-- The tables are generated by the Java application crc32tables in the /java folder
-- LUT2a computes the CRC32s for 64-BIT INPUT WORDS in the form 00 00 00 x 00 00 00 00, where x is the LSB (last received byte)
-- LUT2b computes the CRC32s for 64-BIT INPUT WORDS in the form 00 00 x 00 00 00 00 00 
-- Data bit order: MSb of MSB is first sent/received
-- Note: the returned crc values are NOT inverted and NOT reflected left-right. They are as they would appear
-- when generated by a standard LFSR
---------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity CRC32_LUT2ab is
	 Generic (
		DATA_WIDTH: integer := 32;	
		ADDR_WIDTH: integer := 9
	);
    Port ( 
	    -- Port A
		ADDRA  : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
			-- LUT1a at addresses 0 - 255
			-- LUT1b at addresses 256 - 511
		DOA  : out std_logic_vector(DATA_WIDTH-1 downto 0);

		-- Port B
		ADDRB  : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
			-- LUT1a at addresses 0 - 255
			-- LUT1b at addresses 256 - 511
		DOB  : out std_logic_vector(DATA_WIDTH-1 downto 0)
		);
end entity;

architecture Behavioral of CRC32_LUT2ab is
--------------------------------------------------------
--     SIGNALS
--------------------------------------------------------
-- inferred rom
signal DOA_local: std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
signal DOB_local: std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');
type ROM_TYPE is array ( (2**ADDR_WIDTH)-1 downto 0 ) of std_logic_vector(DATA_WIDTH-1 downto 0);
-- IMPORTANT ORDER INFORMATION: the table below is read from bottom to top and right to left. Thus
-- to restore a common-sense order, address bits are inverted.
constant ROM : ROM_TYPE := (
-- LUT2a
x"00000000", x"490D678D", x"921ACF1A", x"DB17A897", x"20F48383", x"69F9E40E", x"B2EE4C99", x"FBE32B14", 
x"41E90706", x"08E4608B", x"D3F3C81C", x"9AFEAF91", x"611D8485", x"2810E308", x"F3074B9F", x"BA0A2C12", 
x"83D20E0C", x"CADF6981", x"11C8C116", x"58C5A69B", x"A3268D8F", x"EA2BEA02", x"313C4295", x"78312518", 
x"C23B090A", x"8B366E87", x"5021C610", x"192CA19D", x"E2CF8A89", x"ABC2ED04", x"70D54593", x"39D8221E", 
x"036501AF", x"4A686622", x"917FCEB5", x"D872A938", x"2391822C", x"6A9CE5A1", x"B18B4D36", x"F8862ABB", 
x"428C06A9", x"0B816124", x"D096C9B3", x"999BAE3E", x"6278852A", x"2B75E2A7", x"F0624A30", x"B96F2DBD", 
x"80B70FA3", x"C9BA682E", x"12ADC0B9", x"5BA0A734", x"A0438C20", x"E94EEBAD", x"3259433A", x"7B5424B7", 
x"C15E08A5", x"88536F28", x"5344C7BF", x"1A49A032", x"E1AA8B26", x"A8A7ECAB", x"73B0443C", x"3ABD23B1", 
x"06CA035E", x"4FC764D3", x"94D0CC44", x"DDDDABC9", x"263E80DD", x"6F33E750", x"B4244FC7", x"FD29284A", 
x"47230458", x"0E2E63D5", x"D539CB42", x"9C34ACCF", x"67D787DB", x"2EDAE056", x"F5CD48C1", x"BCC02F4C", 
x"85180D52", x"CC156ADF", x"1702C248", x"5E0FA5C5", x"A5EC8ED1", x"ECE1E95C", x"37F641CB", x"7EFB2646", 
x"C4F10A54", x"8DFC6DD9", x"56EBC54E", x"1FE6A2C3", x"E40589D7", x"AD08EE5A", x"761F46CD", x"3F122140", 
x"05AF02F1", x"4CA2657C", x"97B5CDEB", x"DEB8AA66", x"255B8172", x"6C56E6FF", x"B7414E68", x"FE4C29E5", 
x"444605F7", x"0D4B627A", x"D65CCAED", x"9F51AD60", x"64B28674", x"2DBFE1F9", x"F6A8496E", x"BFA52EE3", 
x"867D0CFD", x"CF706B70", x"1467C3E7", x"5D6AA46A", x"A6898F7E", x"EF84E8F3", x"34934064", x"7D9E27E9", 
x"C7940BFB", x"8E996C76", x"558EC4E1", x"1C83A36C", x"E7608878", x"AE6DEFF5", x"757A4762", x"3C7720EF", 
x"0D9406BC", x"44996131", x"9F8EC9A6", x"D683AE2B", x"2D60853F", x"646DE2B2", x"BF7A4A25", x"F6772DA8", 
x"4C7D01BA", x"05706637", x"DE67CEA0", x"976AA92D", x"6C898239", x"2584E5B4", x"FE934D23", x"B79E2AAE", 
x"8E4608B0", x"C74B6F3D", x"1C5CC7AA", x"5551A027", x"AEB28B33", x"E7BFECBE", x"3CA84429", x"75A523A4", 
x"CFAF0FB6", x"86A2683B", x"5DB5C0AC", x"14B8A721", x"EF5B8C35", x"A656EBB8", x"7D41432F", x"344C24A2", 
x"0EF10713", x"47FC609E", x"9CEBC809", x"D5E6AF84", x"2E058490", x"6708E31D", x"BC1F4B8A", x"F5122C07", 
x"4F180015", x"06156798", x"DD02CF0F", x"940FA882", x"6FEC8396", x"26E1E41B", x"FDF64C8C", x"B4FB2B01", 
x"8D23091F", x"C42E6E92", x"1F39C605", x"5634A188", x"ADD78A9C", x"E4DAED11", x"3FCD4586", x"76C0220B", 
x"CCCA0E19", x"85C76994", x"5ED0C103", x"17DDA68E", x"EC3E8D9A", x"A533EA17", x"7E244280", x"3729250D", 
x"0B5E05E2", x"4253626F", x"9944CAF8", x"D049AD75", x"2BAA8661", x"62A7E1EC", x"B9B0497B", x"F0BD2EF6", 
x"4AB702E4", x"03BA6569", x"D8ADCDFE", x"91A0AA73", x"6A438167", x"234EE6EA", x"F8594E7D", x"B15429F0", 
x"888C0BEE", x"C1816C63", x"1A96C4F4", x"539BA379", x"A878886D", x"E175EFE0", x"3A624777", x"736F20FA", 
x"C9650CE8", x"80686B65", x"5B7FC3F2", x"1272A47F", x"E9918F6B", x"A09CE8E6", x"7B8B4071", x"328627FC", 
x"083B044D", x"413663C0", x"9A21CB57", x"D32CACDA", x"28CF87CE", x"61C2E043", x"BAD548D4", x"F3D82F59", 
x"49D2034B", x"00DF64C6", x"DBC8CC51", x"92C5ABDC", x"692680C8", x"202BE745", x"FB3C4FD2", x"B231285F", 
x"8BE90A41", x"C2E46DCC", x"19F3C55B", x"50FEA2D6", x"AB1D89C2", x"E210EE4F", x"390746D8", x"700A2155", 
x"CA000D47", x"830D6ACA", x"581AC25D", x"1117A5D0", x"EAF48EC4", x"A3F9E949", x"78EE41DE", x"31E32653", 
-- LUT2b
x"00000000", x"1B280D78", x"36501AF0", x"2D781788", x"6CA035E0", x"77883898", x"5AF02F10", x"41D82268", 
x"D9406BC0", x"C26866B8", x"EF107130", x"F4387C48", x"B5E05E20", x"AEC85358", x"83B044D0", x"989849A8", 
x"B641CA37", x"AD69C74F", x"8011D0C7", x"9B39DDBF", x"DAE1FFD7", x"C1C9F2AF", x"ECB1E527", x"F799E85F", 
x"6F01A1F7", x"7429AC8F", x"5951BB07", x"4279B67F", x"03A19417", x"1889996F", x"35F18EE7", x"2ED9839F", 
x"684289D9", x"736A84A1", x"5E129329", x"453A9E51", x"04E2BC39", x"1FCAB141", x"32B2A6C9", x"299AABB1", 
x"B102E219", x"AA2AEF61", x"8752F8E9", x"9C7AF591", x"DDA2D7F9", x"C68ADA81", x"EBF2CD09", x"F0DAC071", 
x"DE0343EE", x"C52B4E96", x"E853591E", x"F37B5466", x"B2A3760E", x"A98B7B76", x"84F36CFE", x"9FDB6186", 
x"0743282E", x"1C6B2556", x"311332DE", x"2A3B3FA6", x"6BE31DCE", x"70CB10B6", x"5DB3073E", x"469B0A46", 
x"D08513B2", x"CBAD1ECA", x"E6D50942", x"FDFD043A", x"BC252652", x"A70D2B2A", x"8A753CA2", x"915D31DA", 
x"09C57872", x"12ED750A", x"3F956282", x"24BD6FFA", x"65654D92", x"7E4D40EA", x"53355762", x"481D5A1A", 
x"66C4D985", x"7DECD4FD", x"5094C375", x"4BBCCE0D", x"0A64EC65", x"114CE11D", x"3C34F695", x"271CFBED", 
x"BF84B245", x"A4ACBF3D", x"89D4A8B5", x"92FCA5CD", x"D32487A5", x"C80C8ADD", x"E5749D55", x"FE5C902D", 
x"B8C79A6B", x"A3EF9713", x"8E97809B", x"95BF8DE3", x"D467AF8B", x"CF4FA2F3", x"E237B57B", x"F91FB803", 
x"6187F1AB", x"7AAFFCD3", x"57D7EB5B", x"4CFFE623", x"0D27C44B", x"160FC933", x"3B77DEBB", x"205FD3C3", 
x"0E86505C", x"15AE5D24", x"38D64AAC", x"23FE47D4", x"622665BC", x"790E68C4", x"54767F4C", x"4F5E7234", 
x"D7C63B9C", x"CCEE36E4", x"E196216C", x"FABE2C14", x"BB660E7C", x"A04E0304", x"8D36148C", x"961E19F4", 
x"A5CB3AD3", x"BEE337AB", x"939B2023", x"88B32D5B", x"C96B0F33", x"D243024B", x"FF3B15C3", x"E41318BB", 
x"7C8B5113", x"67A35C6B", x"4ADB4BE3", x"51F3469B", x"102B64F3", x"0B03698B", x"267B7E03", x"3D53737B", 
x"138AF0E4", x"08A2FD9C", x"25DAEA14", x"3EF2E76C", x"7F2AC504", x"6402C87C", x"497ADFF4", x"5252D28C", 
x"CACA9B24", x"D1E2965C", x"FC9A81D4", x"E7B28CAC", x"A66AAEC4", x"BD42A3BC", x"903AB434", x"8B12B94C", 
x"CD89B30A", x"D6A1BE72", x"FBD9A9FA", x"E0F1A482", x"A12986EA", x"BA018B92", x"97799C1A", x"8C519162", 
x"14C9D8CA", x"0FE1D5B2", x"2299C23A", x"39B1CF42", x"7869ED2A", x"6341E052", x"4E39F7DA", x"5511FAA2", 
x"7BC8793D", x"60E07445", x"4D9863CD", x"56B06EB5", x"17684CDD", x"0C4041A5", x"2138562D", x"3A105B55", 
x"A28812FD", x"B9A01F85", x"94D8080D", x"8FF00575", x"CE28271D", x"D5002A65", x"F8783DED", x"E3503095", 
x"754E2961", x"6E662419", x"431E3391", x"58363EE9", x"19EE1C81", x"02C611F9", x"2FBE0671", x"34960B09", 
x"AC0E42A1", x"B7264FD9", x"9A5E5851", x"81765529", x"C0AE7741", x"DB867A39", x"F6FE6DB1", x"EDD660C9", 
x"C30FE356", x"D827EE2E", x"F55FF9A6", x"EE77F4DE", x"AFAFD6B6", x"B487DBCE", x"99FFCC46", x"82D7C13E", 
x"1A4F8896", x"016785EE", x"2C1F9266", x"37379F1E", x"76EFBD76", x"6DC7B00E", x"40BFA786", x"5B97AAFE", 
x"1D0CA0B8", x"0624ADC0", x"2B5CBA48", x"3074B730", x"71AC9558", x"6A849820", x"47FC8FA8", x"5CD482D0", 
x"C44CCB78", x"DF64C600", x"F21CD188", x"E934DCF0", x"A8ECFE98", x"B3C4F3E0", x"9EBCE468", x"8594E910", 
x"AB4D6A8F", x"B06567F7", x"9D1D707F", x"86357D07", x"C7ED5F6F", x"DCC55217", x"F1BD459F", x"EA9548E7", 
x"720D014F", x"69250C37", x"445D1BBF", x"5F7516C7", x"1EAD34AF", x"058539D7", x"28FD2E5F", x"33D52327" 
   	);

--------------------------------------------------------
--      IMPLEMENTATION
--------------------------------------------------------
begin

-- Port A read
DOA <= ROM(to_integer(unsigned(not ADDRA)));	-- see IMPORTANT ORDER INFORMATION above
 

-- Port B read
DOB <= ROM(to_integer(unsigned(not ADDRB)));	-- see IMPORTANT ORDER INFORMATION above

end Behavioral;
